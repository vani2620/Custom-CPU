`ifndef LOGIC_OPERATIONS
`define LOGIC_OPERATIONS
    `define OPCODE_WIDTH    7'h7

    `define ZERO            7'h0
    `define OR              7'h1
    `define AND             7'h2
    `define XOR             7'h3
`endif
