`ifndef ARITHMETIC_OPERATIONS
`define ARITHMETIC_OPERATIONS
    `define OPCODE_WIDTH      7
    `define ADD               7'h08
    `define ADDU              7'h09
    `define SUB               7'h0A
    `define SUBU              7'h0B
    `define MULT              7'h0C
    `define MULTU             7'h0D
    `define DIV               7'h0E
    `define DIVU              7'h0F
`endif
